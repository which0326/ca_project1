module mux1(

);